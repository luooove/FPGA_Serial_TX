module Serial_TEST();

endmodule
